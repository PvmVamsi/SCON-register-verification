package pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	 
         `include "wr_cfg.sv"
         `include "rd_cfg.sv"
         `include "env_cfg.sv"

         `include "wr_xtn.sv"
         `include "wr_mon.sv"
         `include "wr_drv.sv"
         `include "wr_seqr.sv"
         `include "wr_agt.sv"
         `include "wr_agt_top.sv"
         `include "wr_seq.sv"
	
	 `include "rd_xtn.sv"
         `include "rd_mon.sv"
         //`include "rd_driver.sv"
         //`include "rd_seqr.sv"
         `include "rd_agt.sv"
         `include "rd_agt_top.sv"
         //`include "wr_seq.sv"
		
 	 //`include "vseqr.sv"
         //`include "vseq.sv"
         `include "sb.sv"
         `include "env.sv"
	 `include "test.sv"
endpackage
         
	
	  
	 
	 
	
	  
	 
	
	 

